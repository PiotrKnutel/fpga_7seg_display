library verilog;
use verilog.vl_types.all;
entity p06_vlg_vec_tst is
end p06_vlg_vec_tst;
